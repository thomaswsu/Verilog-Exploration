module multipler(input[3:0] X, input[3:0] Y, output[7:0] Z); 
    assign Z = X * Y;
endmodule